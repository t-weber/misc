../../lib/bcd.vhdl