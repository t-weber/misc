../../lib/vga.vhdl