../lib/vga.vhdl