../lib/ram.vhdl