../lib/conv.vhdl