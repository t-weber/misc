../../lib/lfsr.vhdl