../lib/lfsr.vhdl