../lib/clkdiv.vhdl