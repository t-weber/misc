../../lib/ram.vhdl