../../lib/conv.vhdl