../../lib/edge.vhdl