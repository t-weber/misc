../../lib/clkdiv.vhdl