../../lib/sevenseg.vhdl