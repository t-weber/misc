../lib/sevenseg.vhdl