../../lib/div.vhdl