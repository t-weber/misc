../lib/edge.vhdl